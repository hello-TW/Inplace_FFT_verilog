module Inplace_FFT #(
    parameter BW = 16
)(
    input nrst, clk, start, valid,
    input [BW-1:0] inReal, inImag,
    output [BW-1:0]  outReal0, outImag0, outReal1, outImag1
);
    parameter COMP_BW = 2*BW;

    wire we_b0, re_b0, we_b1, re_b1;
    wire [4:0] waddr_b0, waddr_b1, raddr_b0, raddr_b1;
    wire [COMP_BW-1:0] data_in_b0, data_in_b1;
    wire [COMP_BW-1:0] data_out_b0, data_out_b1; 

    simple_dualport_RAM #(COMP_BW) bank0(clk, valid, we_b0, re_b0, waddr_b0, raddr_b0, data_in_b0, data_out_b0);
    simple_dualport_RAM #(COMP_BW) bank1(clk, valid, we_b1, re_b1, waddr_b1, raddr_b1, data_in_b1, data_out_b1);

    Inplace_FFT_core #(BW) core(nrst, clk, start, valid, inReal, inImag, data_out_b0, data_out_b1,
                                we_b0, re_b0, we_b1, re_b1, waddr_b0, waddr_b1, raddr_b0, raddr_b1,
                                data_in_b0, data_in_b1, outReal0, outImag0, outReal1, outImag1);

endmodule
