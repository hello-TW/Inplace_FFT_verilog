library verilog;
use verilog.vl_types.all;
entity Inplace_FFT_tb_sin is
end Inplace_FFT_tb_sin;
